magic
tech sky130A
timestamp 1675880415
<< nwell >>
rect -50 -210 130 -55
<< nmos >>
rect 25 -10 40 50
<< pmos >>
rect 25 -190 40 -80
<< ndiff >>
rect -30 30 25 50
rect -30 10 -25 30
rect -5 10 25 30
rect -30 -10 25 10
rect 40 30 95 50
rect 40 10 70 30
rect 90 10 95 30
rect 40 -10 95 10
<< pdiff >>
rect -30 -130 25 -80
rect -30 -150 -25 -130
rect -5 -150 25 -130
rect -30 -190 25 -150
rect 40 -130 95 -80
rect 40 -150 70 -130
rect 90 -150 95 -130
rect 40 -190 95 -150
<< ndiffc >>
rect -25 10 -5 30
rect 70 10 90 30
<< pdiffc >>
rect -25 -150 -5 -130
rect 70 -150 90 -130
<< poly >>
rect 5 105 60 115
rect 5 70 15 105
rect 50 70 60 105
rect 5 60 60 70
rect 25 50 40 60
rect 25 -80 40 -10
rect 25 -210 40 -190
<< polycont >>
rect 15 70 50 105
<< locali >>
rect 0 105 80 115
rect 0 70 15 105
rect 50 100 165 105
rect 50 80 130 100
rect 150 80 165 100
rect 50 75 165 80
rect 50 70 80 75
rect 0 65 80 70
rect -90 30 5 40
rect -90 10 -85 30
rect -65 10 -25 30
rect -5 10 5 30
rect -90 0 5 10
rect 60 30 110 40
rect 60 10 70 30
rect 90 10 110 30
rect 60 0 110 10
rect 85 -20 110 0
rect 85 -25 120 -20
rect 85 -45 95 -25
rect 115 -45 120 -25
rect 85 -50 120 -45
rect 85 -120 110 -50
rect -90 -130 5 -120
rect -90 -150 -85 -130
rect -65 -150 -25 -130
rect -5 -150 5 -130
rect -90 -160 5 -150
rect 60 -130 110 -120
rect 60 -150 70 -130
rect 90 -150 110 -130
rect 60 -160 110 -150
<< viali >>
rect 130 80 150 100
rect -85 10 -65 30
rect 95 -45 115 -25
rect -85 -150 -65 -130
<< metal1 >>
rect 130 110 150 150
rect 120 100 160 110
rect 120 80 130 100
rect 150 80 160 100
rect 120 70 160 80
rect -110 30 -55 40
rect -110 10 -85 30
rect -65 10 -55 30
rect -110 0 -55 10
rect 85 -20 120 -15
rect 85 -25 185 -20
rect 85 -45 95 -25
rect 115 -45 185 -25
rect 85 -50 185 -45
rect 85 -55 120 -50
rect -115 -130 -50 -120
rect -115 -150 -85 -130
rect -65 -150 -50 -130
rect -115 -160 -50 -150
<< labels >>
rlabel metal1 135 135 145 145 1 in
rlabel metal1 165 -40 175 -30 1 out
rlabel metal1 -110 -145 -100 -135 1 vcc
rlabel metal1 -105 15 -95 25 1 gnd
<< end >>
