Inverter Simulation
* this file edited to remove everything not in tt lib
.lib "/home/kuba/.volare/sky130A/libs.tech/ngspice/sky130.lib.spice" tt

* instantiate the inverter
Xinv OUT IN VGND VPWR VGND INV0

.subckt INV0 out in gnd vcc VSUBS

* NGSPICE file created from mosfet.ext - technology: sky130A


X0 out in gnd VSUBS sky130_fd_pr__nfet_01v8 ad=3.3e+11p pd=2.3e+06u as=3.3e+11p ps=2.3e+06u w=600000u l=150000u
X1 out in vcc w_n100_n420# sky130_fd_pr__pfet_01v8 ad=6.05e+11p pd=3.3e+06u as=6.05e+11p ps=3.3e+06u w=1.1e+06u l=150000u
C0 w_n100_n420# vcc 0.01fF
C1 w_n100_n420# gnd 0.00fF
C2 out vcc 0.02fF
C3 out gnd 0.02fF
C4 w_n100_n420# out 0.02fF
C5 vcc in 0.00fF
C6 gnd in 0.00fF
C7 w_n100_n420# in 0.02fF
C8 out in 0.05fF
C9 gnd vcc 0.05fF
C10 vcc VSUBS 0.12fF
C11 out VSUBS 0.24fF
C12 gnd VSUBS 0.09fF
C13 in VSUBS 0.49fF
C14 w_n100_n420# VSUBS 0.33fF


.ends

* set gnd and power
Vgnd VGND 0 0
Vdd VPWR VGND 1.8

* create pulse
Vin IN VGND pulse(0 1.8 1p 10p 10p 1n 2n)
.tran 10p 2n 0

.control
run
set color0 = white
set color1 = black
plot OUT IN
.endc

.end

