Inverter Simulation
* this file edited to remove everything not in tt lib
.lib "/home/kuba/.volare/sky130A/libs.tech/ngspice/sky130.lib.spice" tt

* instantiate the inverter
Xinv OUT IN VGND VPWR VGND INV0

.subckt INV0 out in gnd vcc VSUBS

